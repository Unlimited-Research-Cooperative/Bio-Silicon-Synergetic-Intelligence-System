library verilog;
use verilog.vl_types.all;
entity generator_vlg_vec_tst is
end generator_vlg_vec_tst;
