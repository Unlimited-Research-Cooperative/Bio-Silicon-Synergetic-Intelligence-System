library verilog;
use verilog.vl_types.all;
entity clock_divider_vlg_vec_tst is
end clock_divider_vlg_vec_tst;
