library verilog;
use verilog.vl_types.all;
entity Parallel_Serial_Converter_vlg_vec_tst is
end Parallel_Serial_Converter_vlg_vec_tst;
