library verilog;
use verilog.vl_types.all;
entity clock_ws_vlg_vec_tst is
end clock_ws_vlg_vec_tst;
